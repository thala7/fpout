------------------------------------------------------------------------------
--  LEON3 Demonstration design
--  Copyright (C) 2013 Aeroflex Gaisler
------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008 - 2014, Aeroflex Gaisler
--  Copyright (C) 2015, Cobham Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;
library techmap;
use techmap.gencomp.all;
use techmap.allclkgen.all;
library gaisler;
use gaisler.memctrl.all;
use gaisler.leon3.all;
use gaisler.uart.all;
use gaisler.misc.all;
use gaisler.spi.all;
use gaisler.net.all;
use gaisler.jtag.all;
--pragma translate_off
use gaisler.sim.all;
--pragma translate_on

library esa;
use esa.memoryctrl.all;
use work.config.all;

entity leon3mp is
  generic (
    fabtech  : integer := CFG_FABTECH;
    memtech  : integer := CFG_MEMTECH;
    padtech  : integer := CFG_PADTECH;
    clktech  : integer := CFG_CLKTECH;
    disas    : integer := CFG_DISAS;     -- Enable disassembly to console
    dbguart  : integer := CFG_DUART;     -- Print UART on console
    pclow    : integer := CFG_PCLOW
    );
  port (
    clk             : in    std_ulogic;
    -- onBoard Cellular RAM, Numonyx StrataFlash and Numonyx Quad Flash
    MemOE           : out   std_ulogic;
    MemWR           : out   std_ulogic;

    RamAdv          : out   std_ulogic;
    RamCS           : out   std_ulogic;
    RamClk          : out   std_ulogic;
    RamCRE          : out   std_ulogic;
    RamLB           : out   std_ulogic;
    RamUB           : out   std_ulogic;
    RamWait         : out   std_ulogic;

    FlashRp         : out   std_ulogic;
    FlashCS         : out   std_ulogic;

    QuadSpiFlashCS  : out   std_ulogic;
    QuadSpiFlashSck : out   std_ulogic;
    QuadSpiFlashDB  : inout std_logic_vector(0 downto 0);

    address         : out   std_logic_vector(25 downto 0);

    data            : inout std_logic_vector(15 downto 0);

    -- 7 segment display
    --seg             : out   std_logic_vector(7 downto 0);
    --an              : out   std_logic_vector(3 downto 0);

    -- LEDs
    led             : out   std_logic_vector(7 downto 0);

    -- Switches
    sw              : in    std_logic_vector(7 downto 0);

    -- Buttons
    btn             : in    std_logic_vector(4 downto 0); -- reset on btn0

    -- VGA Connector
    --vgaRed          : out   std_logic_vector(2 downto 0);
    --vgaGreen        : out   std_logic_vector(2 downto 0);
    --vgaBlue         : out   std_logic_vector(2 downto 1);

    --Hsync           : out   std_ulogic;
    --Vsync           : out   std_ulogic;

    -- 12 pin connectors
    --ja              : inout std_logic_vector(7 downto 0);
    --jb              : inout std_logic_vector(7 downto 0);
    --jc              : inout std_logic_vector(7 downto 0);
    --jd              : inout std_logic_vector(7 downto 0);

    -- SMSC ethernet PHY
    PhyRstn         : out   std_ulogic;
    PhyCrs          : in    std_ulogic;
    PhyCol          : in    std_ulogic;
    PhyClk25Mhz     : out   std_ulogic;

    PhyTxd          : out   std_logic_vector(3 downto 0);
    PhyTxEn         : out   std_ulogic;
    PhyTxClk        : in    std_ulogic;
    PhyTxEr         : out   std_ulogic;

    PhyRxd          : in    std_logic_vector(3 downto 0);
    PhyRxDv         : in    std_ulogic;
    PhyRxEr         : in    std_ulogic;
    PhyRxClk        : in    std_ulogic;

    PhyMdc          : out   std_ulogic;
    PhyMdio         : inout std_logic;


    -- Pic USB-HID interface
    --PS2KeyboardData : inout std_logic;
    --PS2KeyboardClk  : inout std_logic;

    --PS2MouseData    : inout std_logic;
    --PS2MouseClk     : inout std_logic;

    --PicGpio         : out   std_logic_vector(1 downto 0);

    -- USB-RS232 interface
    RsRx            : in    std_logic;
    RsTx            : out   std_logic

    );
end;

architecture rtl of leon3mp is
  signal vcc : std_logic;
  signal gnd : std_logic;

  signal memi : memory_in_type;
  signal memo : memory_out_type;
  signal wpo  : wprot_out_type;

  signal gpioi : gpio_in_type;
  signal gpioo : gpio_out_type;

  signal apbi  : apb_slv_in_type;
  signal apbo  : apb_slv_out_vector := (others => apb_none);
  signal ahbsi : ahb_slv_in_type;
  signal ahbso : ahb_slv_out_vector := (others => ahbs_none);
  signal ahbmi : ahb_mst_in_type;
  signal ahbmo : ahb_mst_out_vector := (others => ahbm_none);

  signal cgi : clkgen_in_type;
  signal cgo : clkgen_out_type;

  signal u1i, dui : uart_in_type;
  signal u1o, duo : uart_out_type;

  signal irqi : irq_in_vector(0 to CFG_NCPU-1);
  signal irqo : irq_out_vector(0 to CFG_NCPU-1);

  signal dbgi : l3_debug_in_vector(0 to CFG_NCPU-1);
  signal dbgo : l3_debug_out_vector(0 to CFG_NCPU-1);

  signal dsui : dsu_in_type;
  signal dsuo : dsu_out_type;

  signal ethi : eth_in_type;
  signal etho : eth_out_type;

  signal gpti : gptimer_in_type;

  signal spii : spi_in_type;
  signal spio : spi_out_type;
  signal slvsel : std_logic_vector(CFG_SPICTRL_SLVS-1 downto 0);

  signal spmi : spimctrl_in_type;
  signal spmo : spimctrl_out_type;

  signal clkm, rstn, clkml  : std_ulogic;
  signal tck, tms, tdi, tdo : std_ulogic;
  signal rstraw             : std_logic;
  signal lock               : std_logic;


-----------start editing-----------------------------
-----------start editing-----------------------------
------------adding tranchecker as component----------
-- component ahbtranschecker is
 -- generic (
    --hindex  : integer := 0;
    --ioaddr  : integer := 16#000#;
    --iomask  : integer := 16#E00#;
    --tech    : integer := DEFMEMTECH; 
    --irq     : integer := 0; 
    --kbytes  : integer := 1); 
  --port (
   -- rst    : in  std_ulogic;
    --clk    : in  std_ulogic;
   -- ahbmi  : in  ahb_mst_in_type;
   --- ahbsi  : in  ahb_slv_in_type;
-------------------------------------------------
    --outccf : out std_logic_vector(31 downto 0);
----------------------------------------------
-------------start editing--------------------
  -- u_tx   : out std_logic;
   --u_tx   : out mini_uart_out_type;
   -- u_rx   : in  std_logic;
    --u_tx   : out std_logic_vector;
   -- u_rx   : in  std_logic_vector;
-------------end editing---------------------
--------------------------------------------
-- ccf_calc_start_port : in std_logic; ----adding this port to make a swicth input
   -- sw_func_or_timed : in std_logic
 -- );
--end component ahbtranschecker;
----------------------------------------
----------end editing------------

-----------------------------------------------------
--component UART_TX is
 -- generic (
  --  g_CLKS_PER_BIT : integer -- := 13920     -- Needs to be set correctly
   -- );
 -- port (
  --  i_Clk       : in  std_logic;
   --- i_TX_DV     : in  std_logic;
--i_TX_Byte   : in  std_logic_vector(7 downto 0);
    --o_TX_Active : out std_logic;
   -- o_TX_Serial : out std_logic;
   -- o_TX_Done   : out std_logic
   --- );
--end component UART_TX;

------------------------------------------------------
----------end editing---------------------------------

  -- RS232 APB Uart
  signal rxd1 : std_logic;
  signal txd1 : std_logic;

-----start editing---
signal outccf_7 : Std_Logic_Vector(31 downto 0); -- Last Byte received--dummy signal
--signal ack_signal : std_logic;---ack signal
--signal IntTx_O_signal : std_logic;---interrupt
--signal Intrx_O_signal : std_logic;---interrupt
--signal WB_DAT_I_SIGNAL: Std_Logic_Vector(7 downto 0); -- Last Byte received
signal ccf_calc_switch_signal : std_logic;--dummy signal
signal sw_func_or_timed : std_logic;--dummy signal

--------------------------------------
----clock divider signals------------
--signal counter : integer :=0;
--signal temp :std_logic :='1'; 
--signal div_clk:std_logic:='1';       
----end editing-----

  
  attribute keep                     : boolean;
  attribute syn_keep                 : boolean;
  attribute syn_preserve             : boolean;
  attribute syn_keep of lock         : signal is true;
  attribute syn_keep of clkml        : signal is true;
  attribute syn_keep of clkm         : signal is true;
  attribute syn_preserve of clkml    : signal is true;
  attribute syn_preserve of clkm     : signal is true;
  attribute keep of lock             : signal is true;
  attribute keep of clkml            : signal is true;
  attribute keep of clkm             : signal is true;

  constant BOARD_FREQ : integer := 100000;                                -- CLK input frequency in KHz
  constant CPU_FREQ   : integer := BOARD_FREQ * CFG_CLKMUL / CFG_CLKDIV;  -- cpu frequency in KHz
begin
--------------------------------------------------------------

----------------------------------------------------------------------
---  Reset and Clock generation  -------------------------------------
----------------------------------------------------------------------

  vcc <= '1';
  gnd <= '0';
---start editing--------------------------------------------
 -- led(7 downto 4) <= (others =>'0'); -- unused leds off
---end editing---------------------------------------------
  
  cgi.pllctrl <= "00";
  cgi.pllrst <= rstraw;

  rst0 : rstgen generic map (acthigh => 1)
    port map (btn(0), clkm, lock, rstn, rstraw);
  lock <= cgo.clklock;
  
  -- clock generator
  clkgen0 : clkgen
    generic map (fabtech, CFG_CLKMUL, CFG_CLKDIV, 0, 0, 0, 0, 0, BOARD_FREQ, 0)
    port map (clk, gnd, clkm, open, open, open, open, cgi, cgo, open, open, open);

---------------------------------------------------------------------- 
---  AHB CONTROLLER --------------------------------------------------
----------------------------------------------------------------------

  ahb0 : ahbctrl
    generic map (defmast => CFG_DEFMST, split => CFG_SPLIT,
                 rrobin  => CFG_RROBIN, ioaddr => CFG_AHBIO, ioen => 1, 
                 nahbm => CFG_NCPU+CFG_AHB_UART+CFG_AHB_JTAG+CFG_GRETH, 
                 nahbs => 8)
    port map (rstn, clkm, ahbmi, ahbmo, ahbsi, ahbso);

----------------------------------------------------------------------
---  LEON3 processor and DSU -----------------------------------------
----------------------------------------------------------------------

  -- LEON3 processor
  leon3gen : if CFG_LEON3 = 1 generate
    cpu : for i in 0 to CFG_NCPU-1 generate
      u0 : leon3s
        generic map (i, fabtech, memtech, CFG_NWIN, CFG_DSU, CFG_FPU, CFG_V8,
                     0, CFG_MAC, pclow, CFG_NOTAG, CFG_NWP, CFG_ICEN, CFG_IREPL, CFG_ISETS, CFG_ILINE,
                     CFG_ISETSZ, CFG_ILOCK, CFG_DCEN, CFG_DREPL, CFG_DSETS, CFG_DLINE, CFG_DSETSZ,
                     CFG_DLOCK, CFG_DSNOOP, CFG_ILRAMEN, CFG_ILRAMSZ, CFG_ILRAMADDR, CFG_DLRAMEN,
                     CFG_DLRAMSZ, CFG_DLRAMADDR, CFG_MMUEN, CFG_ITLBNUM, CFG_DTLBNUM, CFG_TLB_TYPE, CFG_TLB_REP,
                     CFG_LDDEL, disas, CFG_ITBSZ, CFG_PWD, CFG_SVT, CFG_RSTADDR,
                     CFG_NCPU-1, CFG_DFIXED, CFG_SCAN, CFG_MMU_PAGE, CFG_BP, CFG_NP_ASI, CFG_WRPSR)
        port map (clkm, rstn, ahbmi, ahbmo(i), ahbsi, ahbso, irqi(i), irqo(i), dbgi(i), dbgo(i));
    end generate;
---------------------------------------------
---------start editing-----------------------
 --  led(3)  <= not dbgo(0).error;
   -- led(2)  <= not dsuo.active;
---------end editing------------------------
--------------------------------------------

    -- LEON3 Debug Support Unit    
    dsugen : if CFG_DSU = 1 generate
      dsu0 : dsu3
        generic map (hindex => 2, haddr => 16#900#, hmask => 16#F00#,
                     ncpu   => CFG_NCPU, tbits => 30, tech => memtech, irq => 0, kbytes => CFG_ATBSZ)
        port map (rstn, clkm, ahbmi, ahbsi, ahbso(2), dbgo, dbgi, dsui, dsuo);
      dsui.enable <= '1';
    end generate;
  end generate;
  nodsu : if CFG_DSU = 0 generate 
    ahbso(2) <= ahbs_none; dsuo.tstop <= '0'; dsuo.active <= '0';
  end generate;
---------------------------------------------------------------------------------
------------start editing--------------------------------------------------------
   --Debug UART
  dcomgen : if CFG_AHB_UART = 1 generate
    dcom0 : ahbuart
      generic map (hindex => CFG_NCPU, pindex => 4, paddr => 7)
      port map (rstn, clkm, dui, duo, apbi, apbo(4), ahbmi, ahbmo(CFG_NCPU));
    --dsurx_pad : inpad generic map (tech  => padtech) port map (RsRx, dui.rxd);
    --dsutx_pad : outpad generic map (tech => padtech) port map (RsTx, duo.txd);
----------------end editing-------------------------------------------------------
---------------------------------------------
--------start ediitng-----------------------
    --led(0) <= not dui.rxd;
    --led(1) <= not duo.txd;
-------end editing--------------------------
--------------------------------------------
  end generate;
  nouah : if CFG_AHB_UART = 0 generate apbo(4) <= apb_none; end generate;

  ahbjtaggen0 :if CFG_AHB_JTAG = 1 generate
    ahbjtag0 : ahbjtag generic map(tech => fabtech, hindex => CFG_NCPU+CFG_AHB_UART)
      port map(rstn, clkm, tck, tms, tdi, tdo, ahbmi, ahbmo(CFG_NCPU+CFG_AHB_UART),
               open, open, open, open, open, open, open, gnd);
  end generate;

----------------------------------------------------------------------
---  Memory controllers ----------------------------------------------
----------------------------------------------------------------------

  mg2 : if CFG_MCTRL_LEON2 = 1 generate        -- LEON2 memory controller
    sr1 : mctrl generic map (hindex => 5, pindex => 0, paddr => 0, iomask => 0,
        ram8 => CFG_MCTRL_RAM8BIT, ram16 => CFG_MCTRL_RAM16BIT,srbanks=>1)
      port map (rstn, clkm, memi, memo, ahbsi, ahbso(5), apbi, apbo(0), wpo, open);
  end generate;

  memi.brdyn  <= '1';
  memi.bexcn  <= '1';
  memi.writen <= '1';
  memi.wrn    <= "1111";
  memi.bwidth <= "01";

  mg0 : if (CFG_MCTRL_LEON2 = 0) generate 
    apbo(0) <= apb_none;
    ahbso(5) <= ahbs_none;
    memo.bdrive(0) <= '1';
  end generate;

  mgpads : if (CFG_MCTRL_LEON2 /= 0) generate 
    addr_pad : outpadv generic map (tech => padtech, width => 26)
      port map (address, memo.address(26 downto 1));
    oen_pad : outpad generic map (tech => padtech)
      port map (MemOE, memo.oen);
    cs_pad : outpad generic map (tech => padtech)
      port map (RamCS, memo.ramsn(0));
    lb_pad : outpad generic map (tech => padtech)
      port map (RamLB, memo.mben(0));
    ub_pad : outpad generic map (tech => padtech)
      port map (RamUB, memo.mben(1));
    wri_pad : outpad generic map (tech => padtech)
      port map (MemWR, memo.writen);
    fce_pad : outpad generic map (tech => padtech)
      port map (FlashCS, memo.romsn(0));
    frp_pad : outpad generic map (tech => padtech)
      port map (FlashRp, rstn);
  end generate;

  bdr : iopadv generic map (tech => padtech, width => 8)
    port map (data(7 downto 0), memo.data(23 downto 16),
              memo.bdrive(1), memi.data(23 downto 16));
  bdr2 : iopadv generic map (tech => padtech, width => 8)
    port map (data(15 downto 8), memo.data(31 downto 24),
              memo.bdrive(0), memi.data(31 downto 24));
  
  RamCRE <= '0';  
  RamClk <= '0';  
  RamAdv <= '0';



------start editing---------------------------------------------------
-----------start editing-----------------------------
----------------------------------------------------------------------
ahbtc0: entity work.ahbtranschecker
  generic map (
    hindex => 0,
    ioaddr => 16#000#,
    iomask => 16#E00#,
    tech   => CFG_MEMTECH,
    irq    => 0,
    kbytes => 64 )
  port map (
    rst => rstn,
    clk => clkm,
    ahbmi => ahbmi,
    ahbsi =>ahbsi,
    
    outccf => outccf_7,

    u_tx => RsTx,
    ccf_calc_start_port =>ccf_calc_switch_signal,

    sw_func_or_timed => sw_func_or_timed
  );

----------end editing------------

----------------------------------------------------------------------
--miniuart : entity work.UART_TX
  --generic map(
    --g_CLKS_PER_BIT => 870 ---100mhz with 921600br   -- Needs to be set correctly
    --)
  --port map(
    --i_Clk =>clkm,
    --i_TX_DV=>'1',
    --i_TX_Byte =>"01000001",-- DataIn Bus
    --i_TX_Byte =>WB_DAT_I_SIGNAL,-- DataIn Bus
    --o_TX_Active =>IntTx_O_signal ,---dummy signal
    --o_TX_Serial=>RsTx,-- Tx RS232 Line
    --o_TX_Done=>Intrx_O_signal --dummysignal
    --);
---------------------------------------------------------------------
-----------switch for ccf start-----------------------------
    ccf_calc_switch_signal<= sw(7);
--inccf_8_pad : inpadv generic map (tech => padtech, width => 1)
  ---   port map (sw(7), ccf_calc_switch_signal(7));
--------------------------------------------------------------------
 
outccf_8_pad : outpadv generic map (tech => padtech, width => 8)
     port map (led(7 downto 0), outccf_7(7 downto 0));
--------------------------------------------------------------------------------
----------generating continous input---------------------------------
--process(clkm)
 --begin
  --If (clkm'event and clkm='1') then
    -- WB_DAT_I_SIGNAL <= "01000001";
 -- end if;
--end process;

----------------------------------------------------------------------
---------adding clock divider-----------------------------------------
--process (clkm,counter,rstn)
 --begin
 -- if(rstn='0')then counter <=0;temp<='1';
  --  else if(clkm'event and clkm='1')then counter<=counter+1;
    --  if(counter =10000) then temp <= not temp;counter<=0;
      --end if;
  --end if;
 --end if;
 --div_clk<=temp;
--end process;

----------------------------------------------------------------

----------end editing---------------------------------------------------------
    
----------------------------------------------------------------------
---  APB Bridge and various periherals -------------------------------
----------------------------------------------------------------------

  -- APB Bridge
  apb0 : apbctrl
    generic map (hindex => 1, haddr => CFG_APBADDR)
    port map (rstn, clkm, ahbsi, ahbso(1), apbi, apbo);

  -- Interrupt controller
  irqctrl : if CFG_IRQ3_ENABLE /= 0 generate
    irqctrl0 : irqmp
      generic map (pindex => 2, paddr => 2, ncpu => CFG_NCPU)
      port map (rstn, clkm, apbi, apbo(2), irqo, irqi);
  end generate;
  irq3 : if CFG_IRQ3_ENABLE = 0 generate
    x : for i in 0 to CFG_NCPU-1 generate
      irqi(i).irl <= "0000";
    end generate;
    apbo(2) <= apb_none;
  end generate;

  -- Time Unit
  gpt : if CFG_GPT_ENABLE /= 0 generate
    timer0 : gptimer
      generic map (pindex => 3, paddr => 3, pirq => CFG_GPT_IRQ,
                   sepirq => CFG_GPT_SEPIRQ, sbits => CFG_GPT_SW,
                   ntimers => CFG_GPT_NTIM, nbits  => CFG_GPT_TW)
      port map (rstn, clkm, apbi, apbo(3), gpti, open);
    gpti.dhalt  <= dsuo.tstop;
    gpti.extclk <= '0';
  end generate;
  notim : if CFG_GPT_ENABLE = 0 generate apbo(3) <= apb_none; end generate;
---------------------------------------------------------------------------------
----------start editin------------------------------------------------------------

  --Console UART. 
  ua1 : if CFG_UART1_ENABLE /= 0 generate
    uart1 : apbuart                     -- UART 1
      generic map (pindex   => 1, paddr => 1, pirq => 2, console => dbguart, fifosize => CFG_UART1_FIFO)
      port map (rstn, clkm, apbi, apbo(1), u1i, u1o);
    u1i.rxd    <= rxd1;
    u1i.ctsn   <= '0';
    u1i.extclk <= '0';
    txd1       <= u1o.txd;
    -- The USB UART is curently mapped to ahbuart.
   --serrx_pad : inpad generic map (tech  => padtech) port map (RsRx, rxd1);
   --sertx_pad : outpad generic map (tech => padtech) port map (RsTx, txd1);
--   led(0) <= not rxd1;
--    led(1) <= not txd1;
  end generate;
  noua0 : if CFG_UART1_ENABLE = 0 generate apbo(1) <= apb_none; end generate;

  nospi: if CFG_SPICTRL_ENABLE = 0 and CFG_SPIMCTRL = 0 generate
    apbo(7) <= apb_none;
  end generate;

------------------end editing----------------------------------------
-----------------------------------------------------------------------
---  ETHERNET ---------------------------------------------------------
-----------------------------------------------------------------------

  eth0 : if CFG_GRETH = 1 generate -- Gaisler ethernet MAC
    e1 : grethm
      generic map(hindex => CFG_NCPU+CFG_AHB_UART+CFG_AHB_JTAG,
                  pindex => 15, paddr => 15, pirq => 12, memtech => memtech,
                  mdcscaler => CPU_FREQ/1000, enable_mdio => 1, fifosize => CFG_ETH_FIFO,
                  nsync => 1, edcl => CFG_DSU_ETH, edclbufsz => CFG_ETH_BUF,
                  macaddrh => CFG_ETH_ENM, macaddrl => CFG_ETH_ENL, phyrstadr => 7, 
                  ipaddrh => CFG_ETH_IPM, ipaddrl => CFG_ETH_IPL, giga => CFG_GRETH1G)
      port map(rst => rstn, clk => clkm, ahbmi => ahbmi,
               ahbmo => ahbmo(CFG_NCPU+CFG_AHB_UART+CFG_AHB_JTAG), 
               apbi => apbi, apbo => apbo(15), ethi => ethi, etho => etho); 
      PhyRstn<=rstn;
  end generate;

  ethpads : if (CFG_GRETH = 1) generate -- eth pads
    emdio_pad : iopad generic map (tech => padtech)
      port map (PhyMdio, etho.mdio_o, etho.mdio_oe, ethi.mdio_i);
    etxc_pad : clkpad generic map (tech => padtech, arch => 2) 
      port map (PhyTxClk, ethi.tx_clk);
    erxc_pad : clkpad generic map (tech => padtech, arch => 2) 
      port map (PhyRxClk, ethi.rx_clk);
    erxd_pad : inpadv generic map (tech => padtech, width => 4)
      port map (PhyRxd, ethi.rxd(3 downto 0));
    erxdv_pad : inpad generic map (tech => padtech)
      port map (PhyRxDv, ethi.rx_dv);
    erxer_pad : inpad generic map (tech => padtech)
      port map (PhyRxEr, ethi.rx_er);
    erxco_pad : inpad generic map (tech => padtech)
      port map (PhyCol, ethi.rx_col);
    erxcr_pad : inpad generic map (tech => padtech)
      port map (PhyCrs, ethi.rx_crs);

    etxd_pad : outpadv generic map (tech => padtech, width => 4)
      port map (PhyTxd, etho.txd(3 downto 0));
    etxen_pad : outpad generic map (tech => padtech)
      port map (PhyTxEn, etho.tx_en);
    etxer_pad : outpad generic map (tech => padtech)
      port map (PhyTxEr, etho.tx_er);
    emdc_pad : outpad generic map (tech => padtech)
      port map (PhyMdc, etho.mdc);
  end generate;

-----------------------------------------------------------------------
---  AHB ROM ----------------------------------------------------------
-----------------------------------------------------------------------

  bpromgen : if CFG_AHBROMEN /= 0 generate
    brom : entity work.ahbrom
      generic map (hindex => 6, haddr => CFG_AHBRODDR, pipe => CFG_AHBROPIP)
      port map ( rstn, clkm, ahbsi, ahbso(6));
  end generate;
  nobpromgen : if CFG_AHBROMEN = 0 generate
     ahbso(6) <= ahbs_none;
  end generate;

-----------------------------------------------------------------------
---  AHB RAM ----------------------------------------------------------
-----------------------------------------------------------------------

  ahbramgen : if CFG_AHBRAMEN = 1 generate
    ahbram0 : ahbram
      generic map (hindex => 3, haddr => CFG_AHBRADDR, tech => CFG_MEMTECH,
                   kbytes => CFG_AHBRSZ, pipe => CFG_AHBRPIPE)
      port map (rstn, clkm, ahbsi, ahbso(3));
  end generate;
  nram : if CFG_AHBRAMEN = 0 generate ahbso(3) <= ahbs_none; end generate;

-----------------------------------------------------------------------
--  Test report module, only used for simulation ----------------------
-----------------------------------------------------------------------
--pragma translate_off
  test0 : ahbrep generic map (hindex => 4, haddr => 16#200#)
    port map (rstn, clkm, ahbsi, ahbso(4));
--pragma translate_on

-----------------------------------------------------------------------
---  Drive unused bus elements  ---------------------------------------
-----------------------------------------------------------------------

  nam1 : for i in (CFG_NCPU+CFG_AHB_UART+CFG_AHB_JTAG+CFG_GRETH+1) to NAHBMST-1 generate
    ahbmo(i) <= ahbm_none;
  end generate;

-----------------------------------------------------------------------
---  Boot message  ----------------------------------------------------
-----------------------------------------------------------------------

-- pragma translate_off
  x : report_design
    generic map (
      msg1 => "LEON3 Demonstration design for Digilent NEXYS 3 board",
      fabtech => tech_table(fabtech), memtech => tech_table(memtech),
      mdel => 1
      );
-- pragma translate_on

end rtl;
